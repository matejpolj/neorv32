
module vio (
	source);	

	output	[3:0]	source;
endmodule
